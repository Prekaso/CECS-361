
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: CSULB
// Engineers: Jose Aceves & Amin Rezaei
// Create Date: 09/19/2020 06:13:21 PM
// Design Name: 361_Lab3
// Module Name: Lab3
// Revision 0.01 - File Created
//////////////////////////////////////////////////////////////////////////////////


module Lab3(input A, 
            input B,
            input C, 
            input D, 
            input E, 
            output reg Out);
 
    wire S1Ki9SfT3zf2k0NJSnhoYce4t2FloMkXSnhoYce4t2FloMkXK8QYzNIOvoU4vsyuOmeUsdpw8zsRYNyTwj7M3yMfAG1fTClKvgEEfgrolJjhmRsV65zCgyrmxNPUtOFpNg1K2YJUycImgpZvSNwFi0Eh0Px7QUJHWiwSd3owXJPAE6J505IWST2I98nGaqOvuDiixtRkSOMQhLJQaFULkv97biQpAK0MkdASJEUmdEyhTrdmXg1y7b0wxBTEvbeXxrtHmuJFwoxBC4AMyvsPXqmgfGptVwY1TTJQCBBnlwj5G1JSHiYedEWSFRLrhMIhciKBe9OJoFm5r7c4sdlHwBfhkCKb1M6liY92KuXJckLrIUIAhmhIea5jv3OGOs85e3iEcFnxTSQmI671XZp7JIz7HcvLfMl0cFvbzrqBckV6bOpwySJZ0bZMlppD14w1TizSj0PIa07F9mTAeqfo4nJ3kwT2gHcE6wq7VWJsSMRq3lsX7iqTcd0jnGK5gyPwYCjmlCrcgBR9aiX0AecdhgAWYzUZpgFDd7rgE,
    S1Ki9SfT3zf2k0NJSnhoYce4t2FloMkXSnhoYce4t2FloMkXK8QYzNIOvoU4vsyuOmeUsdpw8zsRYNyTwj7M3yMfAG1fTClKvgEEfgrolJjhmRsV65zCgyrmxNPUtOFpNg1K2YJUycImgpZvSNwFi0Eh0Px7QUJHWiwSd3owXJPAE6J505IWST2I98nGaqOvuDiixtRkSOMQhLJQaFULkv97biQpAK0MkdASJEUmdEyhTrdmXg1y7b0wxBTEvbeXxrtHmuJFwoxBC4AMyvsPXqmgfGptVwY1TTJQCBBnlwj5G1JSHiYedEWSFRLrhMIhciKBe9OJoFm5r7c4sdlHwBfhkCKb1M6liY92KuXJckLrIUIAhmhIea5jv3OGOs85e3iEcFnxTSQmI671XZp7JIz7HcvLfMl0cFvbzrqBckV6bOpwySJZ0bZMlppD14wTizSj0PIa07F9mTAeqfo4nJ3kw3T2gHcE6wq7VWJsSMRq3lsX7iqTcd0jnGK5gyPwYCjmlCrcgBR9aiX0AecdhgAWYzUZpgFDd7rgE,
    S1Ki9SfT3zf2k0NJSnhoYce4t2FloMkXSnhoYce4t2FloMkXK8QYzNIOvoU4vsyuOmeUsdpw8zsRYNyTwj7M3yMfAG1fTClKvgEEfgrolJjhmRsV65zCgyrmxNPUtOFpNg1K2YJUycImgpZvSNwFi0Eh0Px7QUJHWiwSd3owXJPAE6J505IWST2I98nGaqOvuDiixtRkSOMQhLJQaFULkv97biQpAK0MkdASJEUmdEyhTrdmXg1y7b0wxBTEvbeXxrtHmuJFwoxBC4AMyvsPXqmgfGptVwY1TTJQCBBnlwj5G1JSHiYedEWSFRLrhMIhciKBe9OJoFm5r7c4sdlHwBfhkCKb1M6liY92KuXJckLrIUIAhmhIea5jv3OGOs85e3iEcFnxTSQmI671XZp7JIz7HcvLfMl0cFvbzrqBckV6bOpwySJZ0bZMlppD14wTizSj0PIa07F9mTAeqfo4nJ3kwT2gHcE6wq7VWJsSMRq3lsX7iqTcd0jnGK5gyPwYCjmlCrcgBR9aiX0AecdhgAWYzUZpgFDpd7rgE,
    S1Ki9SfT3zf2k0NJSnhoYce4t2FloMkXSnhoYce4t2FloMkXK8QYzNIOvoU4vsyuOmeUsdpw8zsRYNyTwj7M3yMfAG1fTClKvgEEfgrolJjhmRsV65zCgyrmxNPUtOFpNg1K2YJUycImgpZvSNwFi0Eh0Px7QUJHWiwSd3owXJPAE6J505IWST2I98nGaqOvuDiixtRkSOMQhLJQaFULkv97biQpAK0MkdASJEUmdEyhTrdmXg1y7b0wxBTEvbeXxrtHmuJFwoxBC4AMyvsPXqmgfGptVwY1TTJQCBBnlwj5G1JSHiYedEWSFRLrhMIhciKBe9OJoFm5r7c4sdlHwBfhkCKb1M6liY92KuXJckLrIUIAhmhIea5jv3OGOs85e3iEcFnxTSQmI671XZp7JIz7HcvLfMl0cFvbzrqBckV6bOpwySJZ0bZMlppD14wTizSj0PIa07F9mTAeqfo4nJ3kwT2gHcE6wq7VWJsSMRq3lsX7iqTcd0jnGK5gyPwYlCjmlCrcgBR9aiX0AecdhgAWYzUZpgFDd7rgE,
    S1Ki9SfT3zf2k0NJSnhoYce4t2FloMkXSnhoYce4t2FloMkXK8QYzNIOvoU4vsyuOmeUsdpw8zsRYNyTwj7M3yMfAG1fTClKvgEEfgrolJjhmRsV65zCgyrmxNPUtOFpNg1K2YJUycImgpZvSNwFi0Eh0Px7QUJHWiwSd3owXJPAE6J505IWST2I98nGaqOvuDiixtRkSOMQhLJQaFULkv97biQpAK0MkdASJEUmdEyhTrdmXg1y7b0wxBTEvbeXxrtHmuJFwoxBC4AMyvsPXqmgfGptVwY1TTJQCBBnlwj5G1JSHiYedEWSFRLrhMIhciKBe9OJoFm5r7c4sdlHwBfhkCKb1M6liY92KuXJckLrIUIAhmhIea5jv3OGOs85e3iEcFnxTSQmI671XZp7JIz7HcvLfMl0cFvbzrqBckV6bOpwySJZ0bZMllppD14wTizSj0PIa07F9mTAeqfo4nJ3kwT2gHcE6wq7VWJsSMRq3lsX7iqTcd0jnGK5gyPwYCjmlCrcgBR9aiX0AecdhgAWYzUZpgFDd7rgE;

    assign S1Ki9SfT3zf2k0NJSnhoYce4t2FloMkXSnhoYce4t2FloMkXK8QYzNIOvoU4vsyuOmeUsdpw8zsRYNyTwj7M3yMfAG1fTClKvgEEfgrolJjhmRsV65zCgyrmxNPUtOFpNg1K2YJUycImgpZvSNwFi0Eh0Px7QUJHWiwSd3owXJPAE6J505IWST2I98nGaqOvuDiixtRkSOMQhLJQaFULkv97biQpAK0MkdASJEUmdEyhTrdmXg1y7b0wxBTEvbeXxrtHmuJFwoxBC4AMyvsPXqmgfGptVwY1TTJQCBBnlwj5G1JSHiYedEWSFRLrhMIhciKBe9OJoFm5r7c4sdlHwBfhkCKb1M6liY92KuXJckLrIUIAhmhIea5jv3OGOs85e3iEcFnxTSQmI671XZp7JIz7HcvLfMl0cFvbzrqBckV6bOpwySJZ0bZMlppD14w1TizSj0PIa07F9mTAeqfo4nJ3kwT2gHcE6wq7VWJsSMRq3lsX7iqTcd0jnGK5gyPwYCjmlCrcgBR9aiX0AecdhgAWYzUZpgFDd7rgE=A;
    assign S1Ki9SfT3zf2k0NJSnhoYce4t2FloMkXSnhoYce4t2FloMkXK8QYzNIOvoU4vsyuOmeUsdpw8zsRYNyTwj7M3yMfAG1fTClKvgEEfgrolJjhmRsV65zCgyrmxNPUtOFpNg1K2YJUycImgpZvSNwFi0Eh0Px7QUJHWiwSd3owXJPAE6J505IWST2I98nGaqOvuDiixtRkSOMQhLJQaFULkv97biQpAK0MkdASJEUmdEyhTrdmXg1y7b0wxBTEvbeXxrtHmuJFwoxBC4AMyvsPXqmgfGptVwY1TTJQCBBnlwj5G1JSHiYedEWSFRLrhMIhciKBe9OJoFm5r7c4sdlHwBfhkCKb1M6liY92KuXJckLrIUIAhmhIea5jv3OGOs85e3iEcFnxTSQmI671XZp7JIz7HcvLfMl0cFvbzrqBckV6bOpwySJZ0bZMlppD14wTizSj0PIa07F9mTAeqfo4nJ3kw3T2gHcE6wq7VWJsSMRq3lsX7iqTcd0jnGK5gyPwYCjmlCrcgBR9aiX0AecdhgAWYzUZpgFDd7rgE=B;
    assign S1Ki9SfT3zf2k0NJSnhoYce4t2FloMkXSnhoYce4t2FloMkXK8QYzNIOvoU4vsyuOmeUsdpw8zsRYNyTwj7M3yMfAG1fTClKvgEEfgrolJjhmRsV65zCgyrmxNPUtOFpNg1K2YJUycImgpZvSNwFi0Eh0Px7QUJHWiwSd3owXJPAE6J505IWST2I98nGaqOvuDiixtRkSOMQhLJQaFULkv97biQpAK0MkdASJEUmdEyhTrdmXg1y7b0wxBTEvbeXxrtHmuJFwoxBC4AMyvsPXqmgfGptVwY1TTJQCBBnlwj5G1JSHiYedEWSFRLrhMIhciKBe9OJoFm5r7c4sdlHwBfhkCKb1M6liY92KuXJckLrIUIAhmhIea5jv3OGOs85e3iEcFnxTSQmI671XZp7JIz7HcvLfMl0cFvbzrqBckV6bOpwySJZ0bZMlppD14wTizSj0PIa07F9mTAeqfo4nJ3kwT2gHcE6wq7VWJsSMRq3lsX7iqTcd0jnGK5gyPwYCjmlCrcgBR9aiX0AecdhgAWYzUZpgFDpd7rgE=C;
    assign S1Ki9SfT3zf2k0NJSnhoYce4t2FloMkXSnhoYce4t2FloMkXK8QYzNIOvoU4vsyuOmeUsdpw8zsRYNyTwj7M3yMfAG1fTClKvgEEfgrolJjhmRsV65zCgyrmxNPUtOFpNg1K2YJUycImgpZvSNwFi0Eh0Px7QUJHWiwSd3owXJPAE6J505IWST2I98nGaqOvuDiixtRkSOMQhLJQaFULkv97biQpAK0MkdASJEUmdEyhTrdmXg1y7b0wxBTEvbeXxrtHmuJFwoxBC4AMyvsPXqmgfGptVwY1TTJQCBBnlwj5G1JSHiYedEWSFRLrhMIhciKBe9OJoFm5r7c4sdlHwBfhkCKb1M6liY92KuXJckLrIUIAhmhIea5jv3OGOs85e3iEcFnxTSQmI671XZp7JIz7HcvLfMl0cFvbzrqBckV6bOpwySJZ0bZMlppD14wTizSj0PIa07F9mTAeqfo4nJ3kwT2gHcE6wq7VWJsSMRq3lsX7iqTcd0jnGK5gyPwYlCjmlCrcgBR9aiX0AecdhgAWYzUZpgFDd7rgE=D;
    assign S1Ki9SfT3zf2k0NJSnhoYce4t2FloMkXSnhoYce4t2FloMkXK8QYzNIOvoU4vsyuOmeUsdpw8zsRYNyTwj7M3yMfAG1fTClKvgEEfgrolJjhmRsV65zCgyrmxNPUtOFpNg1K2YJUycImgpZvSNwFi0Eh0Px7QUJHWiwSd3owXJPAE6J505IWST2I98nGaqOvuDiixtRkSOMQhLJQaFULkv97biQpAK0MkdASJEUmdEyhTrdmXg1y7b0wxBTEvbeXxrtHmuJFwoxBC4AMyvsPXqmgfGptVwY1TTJQCBBnlwj5G1JSHiYedEWSFRLrhMIhciKBe9OJoFm5r7c4sdlHwBfhkCKb1M6liY92KuXJckLrIUIAhmhIea5jv3OGOs85e3iEcFnxTSQmI671XZp7JIz7HcvLfMl0cFvbzrqBckV6bOpwySJZ0bZMllppD14wTizSj0PIa07F9mTAeqfo4nJ3kwT2gHcE6wq7VWJsSMRq3lsX7iqTcd0jnGK5gyPwYCjmlCrcgBR9aiX0AecdhgAWYzUZpgFDd7rgE=E;

    always@(*) begin 
    case({S1Ki9SfT3zf2k0NJSnhoYce4t2FloMkXSnhoYce4t2FloMkXK8QYzNIOvoU4vsyuOmeUsdpw8zsRYNyTwj7M3yMfAG1fTClKvgEEfgrolJjhmRsV65zCgyrmxNPUtOFpNg1K2YJUycImgpZvSNwFi0Eh0Px7QUJHWiwSd3owXJPAE6J505IWST2I98nGaqOvuDiixtRkSOMQhLJQaFULkv97biQpAK0MkdASJEUmdEyhTrdmXg1y7b0wxBTEvbeXxrtHmuJFwoxBC4AMyvsPXqmgfGptVwY1TTJQCBBnlwj5G1JSHiYedEWSFRLrhMIhciKBe9OJoFm5r7c4sdlHwBfhkCKb1M6liY92KuXJckLrIUIAhmhIea5jv3OGOs85e3iEcFnxTSQmI671XZp7JIz7HcvLfMl0cFvbzrqBckV6bOpwySJZ0bZMlppD14wTizSj0PIa07F9mTAeqfo4nJ3kwT2gHcE6wq7VWJsSMRq3lsX7iqTcd0jnGK5gyPwYCjmlCrcgBR9aiX0AecdhgAWYzUZpgFDpd7rgE,
          S1Ki9SfT3zf2k0NJSnhoYce4t2FloMkXSnhoYce4t2FloMkXK8QYzNIOvoU4vsyuOmeUsdpw8zsRYNyTwj7M3yMfAG1fTClKvgEEfgrolJjhmRsV65zCgyrmxNPUtOFpNg1K2YJUycImgpZvSNwFi0Eh0Px7QUJHWiwSd3owXJPAE6J505IWST2I98nGaqOvuDiixtRkSOMQhLJQaFULkv97biQpAK0MkdASJEUmdEyhTrdmXg1y7b0wxBTEvbeXxrtHmuJFwoxBC4AMyvsPXqmgfGptVwY1TTJQCBBnlwj5G1JSHiYedEWSFRLrhMIhciKBe9OJoFm5r7c4sdlHwBfhkCKb1M6liY92KuXJckLrIUIAhmhIea5jv3OGOs85e3iEcFnxTSQmI671XZp7JIz7HcvLfMl0cFvbzrqBckV6bOpwySJZ0bZMlppD14w1TizSj0PIa07F9mTAeqfo4nJ3kwT2gHcE6wq7VWJsSMRq3lsX7iqTcd0jnGK5gyPwYCjmlCrcgBR9aiX0AecdhgAWYzUZpgFDd7rgE,
          S1Ki9SfT3zf2k0NJSnhoYce4t2FloMkXSnhoYce4t2FloMkXK8QYzNIOvoU4vsyuOmeUsdpw8zsRYNyTwj7M3yMfAG1fTClKvgEEfgrolJjhmRsV65zCgyrmxNPUtOFpNg1K2YJUycImgpZvSNwFi0Eh0Px7QUJHWiwSd3owXJPAE6J505IWST2I98nGaqOvuDiixtRkSOMQhLJQaFULkv97biQpAK0MkdASJEUmdEyhTrdmXg1y7b0wxBTEvbeXxrtHmuJFwoxBC4AMyvsPXqmgfGptVwY1TTJQCBBnlwj5G1JSHiYedEWSFRLrhMIhciKBe9OJoFm5r7c4sdlHwBfhkCKb1M6liY92KuXJckLrIUIAhmhIea5jv3OGOs85e3iEcFnxTSQmI671XZp7JIz7HcvLfMl0cFvbzrqBckV6bOpwySJZ0bZMlppD14wTizSj0PIa07F9mTAeqfo4nJ3kw3T2gHcE6wq7VWJsSMRq3lsX7iqTcd0jnGK5gyPwYCjmlCrcgBR9aiX0AecdhgAWYzUZpgFDd7rgE,
          S1Ki9SfT3zf2k0NJSnhoYce4t2FloMkXSnhoYce4t2FloMkXK8QYzNIOvoU4vsyuOmeUsdpw8zsRYNyTwj7M3yMfAG1fTClKvgEEfgrolJjhmRsV65zCgyrmxNPUtOFpNg1K2YJUycImgpZvSNwFi0Eh0Px7QUJHWiwSd3owXJPAE6J505IWST2I98nGaqOvuDiixtRkSOMQhLJQaFULkv97biQpAK0MkdASJEUmdEyhTrdmXg1y7b0wxBTEvbeXxrtHmuJFwoxBC4AMyvsPXqmgfGptVwY1TTJQCBBnlwj5G1JSHiYedEWSFRLrhMIhciKBe9OJoFm5r7c4sdlHwBfhkCKb1M6liY92KuXJckLrIUIAhmhIea5jv3OGOs85e3iEcFnxTSQmI671XZp7JIz7HcvLfMl0cFvbzrqBckV6bOpwySJZ0bZMllppD14wTizSj0PIa07F9mTAeqfo4nJ3kwT2gHcE6wq7VWJsSMRq3lsX7iqTcd0jnGK5gyPwYCjmlCrcgBR9aiX0AecdhgAWYzUZpgFDd7rgE,
          S1Ki9SfT3zf2k0NJSnhoYce4t2FloMkXSnhoYce4t2FloMkXK8QYzNIOvoU4vsyuOmeUsdpw8zsRYNyTwj7M3yMfAG1fTClKvgEEfgrolJjhmRsV65zCgyrmxNPUtOFpNg1K2YJUycImgpZvSNwFi0Eh0Px7QUJHWiwSd3owXJPAE6J505IWST2I98nGaqOvuDiixtRkSOMQhLJQaFULkv97biQpAK0MkdASJEUmdEyhTrdmXg1y7b0wxBTEvbeXxrtHmuJFwoxBC4AMyvsPXqmgfGptVwY1TTJQCBBnlwj5G1JSHiYedEWSFRLrhMIhciKBe9OJoFm5r7c4sdlHwBfhkCKb1M6liY92KuXJckLrIUIAhmhIea5jv3OGOs85e3iEcFnxTSQmI671XZp7JIz7HcvLfMl0cFvbzrqBckV6bOpwySJZ0bZMlppD14wTizSj0PIa07F9mTAeqfo4nJ3kwT2gHcE6wq7VWJsSMRq3lsX7iqTcd0jnGK5gyPwYlCjmlCrcgBR9aiX0AecdhgAWYzUZpgFDd7rgE}) 
          5'b00000 : Out = 1'b1;
          5'b00001 : Out = 1'b1;
          5'b10100 : Out = 1'b1;
          5'b10110 : Out = 1'b1;
          5'b01000 : Out = 1'b1;
          5'b01001 : Out = 1'b1;
          5'b11100 : Out = 1'b1;
          5'b11101 : Out = 1'b1;
          default  : Out = 1'b0;
          endcase
    end
endmodule
